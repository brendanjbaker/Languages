module program;
	initial begin
		$display("Hello, world!");
		$finish;
	end
endmodule
